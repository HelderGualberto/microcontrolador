
--Adder 8 bits
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

ENTITY adder8b is
	port(
		VALUE1    : in  std_logic_vector(7 downto 0);
		VALUE2    : in  std_logic_vector(7 downto 0);
		RESULT	 : out std_logic_vector(7 downto 0);
		OVF : out std_logic := '0'
	);
END;

ARCHITECTURE behavior of adder8b is

signal SUM_AUX, CARRY_AUX: std_logic_vector(7 downto 0);

component FA 
	port 
	   (
			   A, B, C: in std_logic; -- ENTRADAS -> VALOR 1, VALOR 2, CARRY-IN
			   SOMA, CARRY: out std_logic -- SAIDAS -> RESULTADO DA SOMA, CARRY-OUT
			   
		 ); 
end component;

begin
	
	FA1: FA port map (VALUE2(0), VALUE1(0), '0'     , SUM_AUX(0), CARRY_AUX(0));
	FA2: FA port map (VALUE2(1), VALUE1(1), CARRY_AUX(0), SUM_AUX(1), CARRY_AUX(1));
	FA3: FA port map (VALUE2(2), VALUE1(2), CARRY_AUX(1), SUM_AUX(2), CARRY_AUX(2));
	FA4: FA port map (VALUE2(3), VALUE1(3), CARRY_AUX(2), SUM_AUX(3), CARRY_AUX(3));
	FA5: FA port map (VALUE2(4), VALUE1(4), CARRY_AUX(3), SUM_AUX(4), CARRY_AUX(4));
	FA6: FA port map (VALUE2(5), VALUE1(5), CARRY_AUX(4), SUM_AUX(5), CARRY_AUX(5));
	FA7: FA port map (VALUE2(6), VALUE1(6), CARRY_AUX(5), SUM_AUX(6), CARRY_AUX(6));
	FA8: FA port map (VALUE2(7), VALUE1(7), CARRY_AUX(6), SUM_AUX(7), CARRY_AUX(7));
	
	process(CARRY_AUX)
		begin
		
		if (CARRY_AUX(7) = '1') then
			OVF <= '1';
		else
			OVF <= '0';
		END IF;
	end process;
	RESULT <= SUM_AUX;

END behavior;